`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.07.2024 23:37:54
// Design Name: 
// Module Name: Secure_sys_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module secure_sys_tb;
reg [3:0]S,P;
wire GO,STOP;
Secu_Sys uut (.s(S),.p(P),.go(GO),.stop(STOP));
initial
begin
$monitor ("SIMTIME =%g, S=%b,P=%b,GO=%b,STOP=%b", $time,S,P,GO,STOP);
end
initial begin
#5 S =4'b0000; P=4'b0000;
#5 S =4'b0000; P=4'b0001;
#5 S =4'b0000; P=4'b0010;
#5 S =4'b0000; P=4'b0011;
#5 S =4'b0000; P=4'b0100;
#5 S =4'b0000; P=4'b0101;
#5 S =4'b0000; P=4'b0110;
#5 S =4'b0000; P=4'b0111;
#5 S =4'b0000; P=4'b1000;
#5 S =4'b0000; P=4'b1001;
#5 S =4'b0000; P=4'b1010;
#5 S =4'b0000; P=4'b1011;
#5 S =4'b0000; P=4'b1100;
#5 S =4'b0000; P=4'b1101;
#5 S =4'b0000; P=4'b1110;
#5 S =4'b0000; P=4'b1111;


#5 S =4'b0001; P=4'b0000;
#5 S =4'b0001; P=4'b0001;
#5 S =4'b0001; P=4'b0010;
#5 S =4'b0001; P=4'b0011;
#5 S =4'b0001; P=4'b0100;
#5 S =4'b0001; P=4'b0101;
#5 S =4'b0001; P=4'b0110;
#5 S =4'b0001; P=4'b0111;
#5 S =4'b0001; P=4'b1000;
#5 S =4'b0001; P=4'b1001;
#5 S =4'b0001; P=4'b1010;
#5 S =4'b0001; P=4'b1011;
#5 S =4'b0001; P=4'b1100;
#5 S =4'b0001; P=4'b1101;
#5 S =4'b0001; P=4'b1110;
#5 S =4'b0001; P=4'b1111;

#5 S =4'b0010; P=4'b0000;
#5 S =4'b0010; P=4'b0001;
#5 S =4'b0010; P=4'b0010;
#5 S =4'b0010; P=4'b0011;
#5 S =4'b0010; P=4'b0100;
#5 S =4'b0010; P=4'b0101;
#5 S =4'b0010; P=4'b0110;
#5 S =4'b0010; P=4'b0111;
#5 S =4'b0010; P=4'b1000;
#5 S =4'b0010; P=4'b1001;
#5 S =4'b0010; P=4'b1010;
#5 S =4'b0010; P=4'b1011;
#5 S =4'b0010; P=4'b1100;
#5 S =4'b0010; P=4'b1101;
#5 S =4'b0010; P=4'b1110;
#5 S =4'b0010; P=4'b1111;

#5 S =4'b0011; P=4'b0000;
#5 S =4'b0011; P=4'b0001;
#5 S =4'b0011; P=4'b0010;
#5 S =4'b0011; P=4'b0011;
#5 S =4'b0011; P=4'b0100;
#5 S =4'b0011; P=4'b0101;
#5 S =4'b0011; P=4'b0110;
#5 S =4'b0011; P=4'b0111;
#5 S =4'b0011; P=4'b1000;
#5 S =4'b0011; P=4'b1001;
#5 S =4'b0011; P=4'b1010;
#5 S =4'b0011; P=4'b1011;
#5 S =4'b0011; P=4'b1100;
#5 S =4'b0011; P=4'b1101;
#5 S =4'b0011; P=4'b1110;
#5 S =4'b0011; P=4'b1111;

#5 S =4'b0100; P=4'b0000;
#5 S =4'b0100; P=4'b0001;
#5 S =4'b0100; P=4'b0010;
#5 S =4'b0100; P=4'b0011;
#5 S =4'b0100; P=4'b0100;
#5 S =4'b0100; P=4'b0101;
#5 S =4'b0100; P=4'b0110;
#5 S =4'b0100; P=4'b0111;
#5 S =4'b0100; P=4'b1000;
#5 S =4'b0100; P=4'b1001;
#5 S =4'b0100; P=4'b1010;
#5 S =4'b0100; P=4'b1011;
#5 S =4'b0100; P=4'b1100;
#5 S =4'b0100; P=4'b1101;
#5 S =4'b0100; P=4'b1110;
#5 S =4'b0100; P=4'b1111;

#5 S =4'b0101; P=4'b0000;
#5 S =4'b0101; P=4'b0001;
#5 S =4'b0101; P=4'b0010;
#5 S =4'b0101; P=4'b0011;
#5 S =4'b0101; P=4'b0100;
#5 S =4'b0101; P=4'b0101;
#5 S =4'b0101; P=4'b0110;
#5 S =4'b0101; P=4'b0111;
#5 S =4'b0101; P=4'b1000;
#5 S =4'b0101; P=4'b1001;
#5 S =4'b0101; P=4'b1010;
#5 S =4'b0101; P=4'b1011;
#5 S =4'b0101; P=4'b1100;
#5 S =4'b0101; P=4'b1101;
#5 S =4'b0101; P=4'b1110;
#5 S =4'b0101; P=4'b1111;

#5 S =4'b0110; P=4'b0000;
#5 S =4'b0110; P=4'b0001;
#5 S =4'b0110; P=4'b0010;
#5 S =4'b0110; P=4'b0011;
#5 S =4'b0110; P=4'b0100;
#5 S =4'b0110; P=4'b0101;
#5 S =4'b0110; P=4'b0110;
#5 S =4'b0110; P=4'b0111;
#5 S =4'b0110; P=4'b1000;
#5 S =4'b0110; P=4'b1001;
#5 S =4'b0110; P=4'b1010;
#5 S =4'b0110; P=4'b1011;
#5 S =4'b0110; P=4'b1100;
#5 S =4'b0110; P=4'b1101;
#5 S =4'b0110; P=4'b1110;
#5 S =4'b0110; P=4'b1111;

#5 S =4'b0111; P=4'b0000;
#5 S =4'b0111; P=4'b0001;
#5 S =4'b0111; P=4'b0010;
#5 S =4'b0111; P=4'b0011;
#5 S =4'b0111; P=4'b0100;
#5 S =4'b0111; P=4'b0101;
#5 S =4'b0111; P=4'b0110;
#5 S =4'b0111; P=4'b0111;
#5 S =4'b0111; P=4'b1000;
#5 S =4'b0111; P=4'b1001;
#5 S =4'b0111; P=4'b1010;
#5 S =4'b0111; P=4'b1011;
#5 S =4'b0111; P=4'b1100;
#5 S =4'b0111; P=4'b1101;
#5 S =4'b0111; P=4'b1110;
#5 S =4'b0111; P=4'b1111;

#5 S =4'b1000; P=4'b0000;
#5 S =4'b1000; P=4'b0001;
#5 S =4'b1000; P=4'b0010;
#5 S =4'b1000; P=4'b0011;
#5 S =4'b1000; P=4'b0100;
#5 S =4'b1000; P=4'b0101;
#5 S =4'b1000; P=4'b0110;
#5 S =4'b1000; P=4'b0111;
#5 S =4'b1000; P=4'b1000;
#5 S =4'b1000; P=4'b1001;
#5 S =4'b1000; P=4'b1010;
#5 S =4'b1000; P=4'b1011;
#5 S =4'b1000; P=4'b1100;
#5 S =4'b1000; P=4'b1101;
#5 S =4'b1000; P=4'b1110;
#5 S =4'b1000; P=4'b1111;

#5 S =4'b1001; P=4'b0000;
#5 S =4'b1001; P=4'b0001;
#5 S =4'b1001; P=4'b0010;
#5 S =4'b1001; P=4'b0011;
#5 S =4'b1001; P=4'b0100;
#5 S =4'b1001; P=4'b0101;
#5 S =4'b1001; P=4'b0110;
#5 S =4'b1001; P=4'b0111;
#5 S =4'b1001; P=4'b1000;
#5 S =4'b1001; P=4'b1001;
#5 S =4'b1001; P=4'b1010;
#5 S =4'b1001; P=4'b1011;
#5 S =4'b1001; P=4'b1100;
#5 S =4'b1001; P=4'b1101;
#5 S =4'b1001; P=4'b1110;
#5 S =4'b1001; P=4'b1111;

#5 S =4'b1010; P=4'b0000;
#5 S =4'b1010; P=4'b0001;
#5 S =4'b1010; P=4'b0010;
#5 S =4'b1010; P=4'b0011;
#5 S =4'b1010; P=4'b0100;
#5 S =4'b1010; P=4'b0101;
#5 S =4'b1010; P=4'b0110;
#5 S =4'b1010; P=4'b0111;
#5 S =4'b1010; P=4'b1000;
#5 S =4'b1010; P=4'b1001;
#5 S =4'b1010; P=4'b1010;
#5 S =4'b1010; P=4'b1011;
#5 S =4'b1010; P=4'b1100;
#5 S =4'b1010; P=4'b1101;
#5 S =4'b1010; P=4'b1110;
#5 S =4'b1010; P=4'b1111;

#5 S =4'b1011; P=4'b0000;
#5 S =4'b1011; P=4'b0001;
#5 S =4'b1011; P=4'b0010;
#5 S =4'b1011; P=4'b0011;
#5 S =4'b1011; P=4'b0100;
#5 S =4'b1011; P=4'b0101;
#5 S =4'b1011; P=4'b0110;
#5 S =4'b1011; P=4'b0111;
#5 S =4'b1011; P=4'b1000;
#5 S =4'b1011; P=4'b1001;
#5 S =4'b1011; P=4'b1010;
#5 S =4'b1011; P=4'b1011;
#5 S =4'b1011; P=4'b1100;
#5 S =4'b1011; P=4'b1101;
#5 S =4'b1011; P=4'b1110;
#5 S =4'b1011; P=4'b1111;

#5 S =4'b1100; P=4'b0000;
#5 S =4'b1100; P=4'b0001;
#5 S =4'b1100; P=4'b0010;
#5 S =4'b1100; P=4'b0011;
#5 S =4'b1100; P=4'b0100;
#5 S =4'b1100; P=4'b0101;
#5 S =4'b1100; P=4'b0110;
#5 S =4'b1100; P=4'b0111;
#5 S =4'b1100; P=4'b1000;
#5 S =4'b1100; P=4'b1001;
#5 S =4'b1100; P=4'b1010;
#5 S =4'b1100; P=4'b1011;
#5 S =4'b1100; P=4'b1100;
#5 S =4'b1100; P=4'b1101;
#5 S =4'b1100; P=4'b1110;
#5 S =4'b1100; P=4'b1111;

#5 S =4'b1101; P=4'b0000;
#5 S =4'b1101; P=4'b0001;
#5 S =4'b1101; P=4'b0010;
#5 S =4'b1101; P=4'b0011;
#5 S =4'b1101; P=4'b0100;
#5 S =4'b1101; P=4'b0101;
#5 S =4'b1101; P=4'b0110;
#5 S =4'b1101; P=4'b0111;
#5 S =4'b1101; P=4'b1000;
#5 S =4'b1101; P=4'b1001;
#5 S =4'b1101; P=4'b1010;
#5 S =4'b1101; P=4'b1011;
#5 S =4'b1101; P=4'b1100;
#5 S =4'b1101; P=4'b1101;
#5 S =4'b1101; P=4'b1110;
#5 S =4'b1101; P=4'b1111;

#5 S =4'b1110; P=4'b0000;
#5 S =4'b1110; P=4'b0001;
#5 S =4'b1110; P=4'b0010;
#5 S =4'b1110; P=4'b0011;
#5 S =4'b1110; P=4'b0100;
#5 S =4'b1110; P=4'b0101;
#5 S =4'b1110; P=4'b0110;
#5 S =4'b1110; P=4'b0111;
#5 S =4'b1110; P=4'b1000;
#5 S =4'b1110; P=4'b1001;
#5 S =4'b1110; P=4'b1010;
#5 S =4'b1110; P=4'b1011;
#5 S =4'b1110; P=4'b1100;
#5 S =4'b1110; P=4'b1101;
#5 S =4'b1110; P=4'b1110;
#5 S =4'b1110; P=4'b1111;

#5 S =4'b1111; P=4'b0000;
#5 S =4'b1111; P=4'b0001;
#5 S =4'b1111; P=4'b0010;
#5 S =4'b1111; P=4'b0011;
#5 S =4'b1111; P=4'b0100;
#5 S =4'b1111; P=4'b0101;
#5 S =4'b1111; P=4'b0110;
#5 S =4'b1111; P=4'b0111;
#5 S =4'b1111; P=4'b1000;
#5 S =4'b1111; P=4'b1001;
#5 S =4'b1111; P=4'b1010;
#5 S =4'b1111; P=4'b1011;
#5 S =4'b1111; P=4'b1100;
#5 S =4'b1111; P=4'b1101;
#5 S =4'b1111; P=4'b1110;
#5 S =4'b1111; P=4'b1111;

end 
endmodule

